module test(input logic test);
	always test before use;
endmodule